package lwdo_regs_rtl_pkg;
  localparam int SYS_MAGIC_BYTE_WIDTH = 4;
  localparam int SYS_MAGIC_BYTE_SIZE = 4;
  localparam bit [8:0] SYS_MAGIC_BYTE_OFFSET = 9'h000;
  localparam int SYS_MAGIC_MAGIC_BIT_WIDTH = 32;
  localparam bit [31:0] SYS_MAGIC_MAGIC_BIT_MASK = 32'hffffffff;
  localparam int SYS_MAGIC_MAGIC_BIT_OFFSET = 0;
  localparam int SYS_VERSION_BYTE_WIDTH = 4;
  localparam int SYS_VERSION_BYTE_SIZE = 4;
  localparam bit [8:0] SYS_VERSION_BYTE_OFFSET = 9'h004;
  localparam int SYS_VERSION_MAJOR_BIT_WIDTH = 16;
  localparam bit [15:0] SYS_VERSION_MAJOR_BIT_MASK = 16'hffff;
  localparam int SYS_VERSION_MAJOR_BIT_OFFSET = 0;
  localparam int SYS_VERSION_MINOR_BIT_WIDTH = 16;
  localparam bit [15:0] SYS_VERSION_MINOR_BIT_MASK = 16'hffff;
  localparam int SYS_VERSION_MINOR_BIT_OFFSET = 16;
  localparam int SYS_CON_BYTE_WIDTH = 2;
  localparam int SYS_CON_BYTE_SIZE = 2;
  localparam bit [8:0] SYS_CON_BYTE_OFFSET = 9'h008;
  localparam int SYS_CON_SYS_RST_BIT_WIDTH = 1;
  localparam bit SYS_CON_SYS_RST_BIT_MASK = 1'h1;
  localparam int SYS_CON_SYS_RST_BIT_OFFSET = 0;
  localparam int SYS_PLL_BYTE_WIDTH = 2;
  localparam int SYS_PLL_BYTE_SIZE = 2;
  localparam bit [8:0] SYS_PLL_BYTE_OFFSET = 9'h00a;
  localparam int SYS_PLL_DIVR_BIT_WIDTH = 4;
  localparam bit [3:0] SYS_PLL_DIVR_BIT_MASK = 4'hf;
  localparam int SYS_PLL_DIVR_BIT_OFFSET = 0;
  localparam int SYS_PLL_DIVF_BIT_WIDTH = 7;
  localparam bit [6:0] SYS_PLL_DIVF_BIT_MASK = 7'h7f;
  localparam int SYS_PLL_DIVF_BIT_OFFSET = 4;
  localparam int SYS_PLL_DIVQ_BIT_WIDTH = 3;
  localparam bit [2:0] SYS_PLL_DIVQ_BIT_MASK = 3'h7;
  localparam int SYS_PLL_DIVQ_BIT_OFFSET = 11;
  localparam int PDET_CON_BYTE_WIDTH = 2;
  localparam int PDET_CON_BYTE_SIZE = 2;
  localparam bit [8:0] PDET_CON_BYTE_OFFSET = 9'h020;
  localparam int PDET_CON_EN_BIT_WIDTH = 1;
  localparam bit PDET_CON_EN_BIT_MASK = 1'h1;
  localparam int PDET_CON_EN_BIT_OFFSET = 0;
  localparam int PDET_CON_ECLK2_SLOW_BIT_WIDTH = 1;
  localparam bit PDET_CON_ECLK2_SLOW_BIT_MASK = 1'h1;
  localparam int PDET_CON_ECLK2_SLOW_BIT_OFFSET = 1;
  localparam int PDET_N1_BYTE_WIDTH = 4;
  localparam int PDET_N1_BYTE_SIZE = 4;
  localparam bit [8:0] PDET_N1_BYTE_OFFSET = 9'h022;
  localparam int PDET_N1_VAL_BIT_WIDTH = 32;
  localparam bit [31:0] PDET_N1_VAL_BIT_MASK = 32'hffffffff;
  localparam int PDET_N1_VAL_BIT_OFFSET = 0;
  localparam int PDET_N2_BYTE_WIDTH = 4;
  localparam int PDET_N2_BYTE_SIZE = 4;
  localparam bit [8:0] PDET_N2_BYTE_OFFSET = 9'h026;
  localparam int PDET_N2_VAL_BIT_WIDTH = 32;
  localparam bit [31:0] PDET_N2_VAL_BIT_MASK = 32'hffffffff;
  localparam int PDET_N2_VAL_BIT_OFFSET = 0;
  localparam int ADCT_CON_BYTE_WIDTH = 2;
  localparam int ADCT_CON_BYTE_SIZE = 2;
  localparam bit [8:0] ADCT_CON_BYTE_OFFSET = 9'h040;
  localparam int ADCT_CON_SRATE1_EN_BIT_WIDTH = 1;
  localparam bit ADCT_CON_SRATE1_EN_BIT_MASK = 1'h1;
  localparam int ADCT_CON_SRATE1_EN_BIT_OFFSET = 0;
  localparam int ADCT_CON_SRATE2_EN_BIT_WIDTH = 1;
  localparam bit ADCT_CON_SRATE2_EN_BIT_MASK = 1'h1;
  localparam int ADCT_CON_SRATE2_EN_BIT_OFFSET = 1;
  localparam int ADCT_CON_PULS1_EN_BIT_WIDTH = 1;
  localparam bit ADCT_CON_PULS1_EN_BIT_MASK = 1'h1;
  localparam int ADCT_CON_PULS1_EN_BIT_OFFSET = 2;
  localparam int ADCT_CON_PULS2_EN_BIT_WIDTH = 1;
  localparam bit ADCT_CON_PULS2_EN_BIT_MASK = 1'h1;
  localparam int ADCT_CON_PULS2_EN_BIT_OFFSET = 3;
  localparam int ADCT_SRATE1_PSC_DIV_BYTE_WIDTH = 2;
  localparam int ADCT_SRATE1_PSC_DIV_BYTE_SIZE = 2;
  localparam bit [8:0] ADCT_SRATE1_PSC_DIV_BYTE_OFFSET = 9'h042;
  localparam int ADCT_SRATE1_PSC_DIV_VAL_BIT_WIDTH = 8;
  localparam bit [7:0] ADCT_SRATE1_PSC_DIV_VAL_BIT_MASK = 8'hff;
  localparam int ADCT_SRATE1_PSC_DIV_VAL_BIT_OFFSET = 0;
  localparam int ADCT_SRATE2_PSC_DIV_BYTE_WIDTH = 2;
  localparam int ADCT_SRATE2_PSC_DIV_BYTE_SIZE = 2;
  localparam bit [8:0] ADCT_SRATE2_PSC_DIV_BYTE_OFFSET = 9'h044;
  localparam int ADCT_SRATE2_PSC_DIV_VAL_BIT_WIDTH = 8;
  localparam bit [7:0] ADCT_SRATE2_PSC_DIV_VAL_BIT_MASK = 8'hff;
  localparam int ADCT_SRATE2_PSC_DIV_VAL_BIT_OFFSET = 0;
  localparam int ADCT_PULS1_PSC_DIV_BYTE_WIDTH = 4;
  localparam int ADCT_PULS1_PSC_DIV_BYTE_SIZE = 4;
  localparam bit [8:0] ADCT_PULS1_PSC_DIV_BYTE_OFFSET = 9'h046;
  localparam int ADCT_PULS1_PSC_DIV_VAL_BIT_WIDTH = 23;
  localparam bit [22:0] ADCT_PULS1_PSC_DIV_VAL_BIT_MASK = 23'h7fffff;
  localparam int ADCT_PULS1_PSC_DIV_VAL_BIT_OFFSET = 0;
  localparam int ADCT_PULS2_PSC_DIV_BYTE_WIDTH = 4;
  localparam int ADCT_PULS2_PSC_DIV_BYTE_SIZE = 4;
  localparam bit [8:0] ADCT_PULS2_PSC_DIV_BYTE_OFFSET = 9'h04a;
  localparam int ADCT_PULS2_PSC_DIV_VAL_BIT_WIDTH = 23;
  localparam bit [22:0] ADCT_PULS2_PSC_DIV_VAL_BIT_MASK = 23'h7fffff;
  localparam int ADCT_PULS2_PSC_DIV_VAL_BIT_OFFSET = 0;
  localparam int ADCT_PULS1_DLY_BYTE_WIDTH = 2;
  localparam int ADCT_PULS1_DLY_BYTE_SIZE = 2;
  localparam bit [8:0] ADCT_PULS1_DLY_BYTE_OFFSET = 9'h04e;
  localparam int ADCT_PULS1_DLY_VAL_BIT_WIDTH = 9;
  localparam bit [8:0] ADCT_PULS1_DLY_VAL_BIT_MASK = 9'h1ff;
  localparam int ADCT_PULS1_DLY_VAL_BIT_OFFSET = 0;
  localparam int ADCT_PULS2_DLY_BYTE_WIDTH = 2;
  localparam int ADCT_PULS2_DLY_BYTE_SIZE = 2;
  localparam bit [8:0] ADCT_PULS2_DLY_BYTE_OFFSET = 9'h050;
  localparam int ADCT_PULS2_DLY_VAL_BIT_WIDTH = 9;
  localparam bit [8:0] ADCT_PULS2_DLY_VAL_BIT_MASK = 9'h1ff;
  localparam int ADCT_PULS2_DLY_VAL_BIT_OFFSET = 0;
  localparam int ADCT_PULS1_PWIDTH_BYTE_WIDTH = 2;
  localparam int ADCT_PULS1_PWIDTH_BYTE_SIZE = 2;
  localparam bit [8:0] ADCT_PULS1_PWIDTH_BYTE_OFFSET = 9'h052;
  localparam int ADCT_PULS1_PWIDTH_VAL_BIT_WIDTH = 16;
  localparam bit [15:0] ADCT_PULS1_PWIDTH_VAL_BIT_MASK = 16'hffff;
  localparam int ADCT_PULS1_PWIDTH_VAL_BIT_OFFSET = 0;
  localparam int ADCT_PULS2_PWIDTH_BYTE_WIDTH = 2;
  localparam int ADCT_PULS2_PWIDTH_BYTE_SIZE = 2;
  localparam bit [8:0] ADCT_PULS2_PWIDTH_BYTE_OFFSET = 9'h054;
  localparam int ADCT_PULS2_PWIDTH_VAL_BIT_WIDTH = 16;
  localparam bit [15:0] ADCT_PULS2_PWIDTH_VAL_BIT_MASK = 16'hffff;
  localparam int ADCT_PULS2_PWIDTH_VAL_BIT_OFFSET = 0;
  localparam int ADC_CON_BYTE_WIDTH = 2;
  localparam int ADC_CON_BYTE_SIZE = 2;
  localparam bit [8:0] ADC_CON_BYTE_OFFSET = 9'h080;
  localparam int ADC_CON_ADC1_EN_BIT_WIDTH = 1;
  localparam bit ADC_CON_ADC1_EN_BIT_MASK = 1'h1;
  localparam int ADC_CON_ADC1_EN_BIT_OFFSET = 0;
  localparam int ADC_CON_ADC2_EN_BIT_WIDTH = 1;
  localparam bit ADC_CON_ADC2_EN_BIT_MASK = 1'h1;
  localparam int ADC_CON_ADC2_EN_BIT_OFFSET = 1;
  localparam int ADC_FIFO1_STS_BYTE_WIDTH = 2;
  localparam int ADC_FIFO1_STS_BYTE_SIZE = 2;
  localparam bit [8:0] ADC_FIFO1_STS_BYTE_OFFSET = 9'h082;
  localparam int ADC_FIFO1_STS_EMPTY_BIT_WIDTH = 1;
  localparam bit ADC_FIFO1_STS_EMPTY_BIT_MASK = 1'h1;
  localparam int ADC_FIFO1_STS_EMPTY_BIT_OFFSET = 0;
  localparam int ADC_FIFO1_STS_FULL_BIT_WIDTH = 1;
  localparam bit ADC_FIFO1_STS_FULL_BIT_MASK = 1'h1;
  localparam int ADC_FIFO1_STS_FULL_BIT_OFFSET = 1;
  localparam int ADC_FIFO1_STS_HFULL_BIT_WIDTH = 1;
  localparam bit ADC_FIFO1_STS_HFULL_BIT_MASK = 1'h1;
  localparam int ADC_FIFO1_STS_HFULL_BIT_OFFSET = 2;
  localparam int ADC_FIFO1_STS_OVFL_BIT_WIDTH = 1;
  localparam bit ADC_FIFO1_STS_OVFL_BIT_MASK = 1'h1;
  localparam int ADC_FIFO1_STS_OVFL_BIT_OFFSET = 3;
  localparam int ADC_FIFO1_STS_UDFL_BIT_WIDTH = 1;
  localparam bit ADC_FIFO1_STS_UDFL_BIT_MASK = 1'h1;
  localparam int ADC_FIFO1_STS_UDFL_BIT_OFFSET = 4;
  localparam int ADC_FIFO2_STS_BYTE_WIDTH = 2;
  localparam int ADC_FIFO2_STS_BYTE_SIZE = 2;
  localparam bit [8:0] ADC_FIFO2_STS_BYTE_OFFSET = 9'h084;
  localparam int ADC_FIFO2_STS_EMPTY_BIT_WIDTH = 1;
  localparam bit ADC_FIFO2_STS_EMPTY_BIT_MASK = 1'h1;
  localparam int ADC_FIFO2_STS_EMPTY_BIT_OFFSET = 0;
  localparam int ADC_FIFO2_STS_FULL_BIT_WIDTH = 1;
  localparam bit ADC_FIFO2_STS_FULL_BIT_MASK = 1'h1;
  localparam int ADC_FIFO2_STS_FULL_BIT_OFFSET = 1;
  localparam int ADC_FIFO2_STS_HFULL_BIT_WIDTH = 1;
  localparam bit ADC_FIFO2_STS_HFULL_BIT_MASK = 1'h1;
  localparam int ADC_FIFO2_STS_HFULL_BIT_OFFSET = 2;
  localparam int ADC_FIFO2_STS_OVFL_BIT_WIDTH = 1;
  localparam bit ADC_FIFO2_STS_OVFL_BIT_MASK = 1'h1;
  localparam int ADC_FIFO2_STS_OVFL_BIT_OFFSET = 3;
  localparam int ADC_FIFO2_STS_UDFL_BIT_WIDTH = 1;
  localparam bit ADC_FIFO2_STS_UDFL_BIT_MASK = 1'h1;
  localparam int ADC_FIFO2_STS_UDFL_BIT_OFFSET = 4;
  localparam int FTUN_VTUNE_SET_BYTE_WIDTH = 2;
  localparam int FTUN_VTUNE_SET_BYTE_SIZE = 2;
  localparam bit [8:0] FTUN_VTUNE_SET_BYTE_OFFSET = 9'h0a0;
  localparam int FTUN_VTUNE_SET_VAL_BIT_WIDTH = 16;
  localparam bit [15:0] FTUN_VTUNE_SET_VAL_BIT_MASK = 16'hffff;
  localparam int FTUN_VTUNE_SET_VAL_BIT_OFFSET = 0;
  localparam int TEST_RW1_BYTE_WIDTH = 2;
  localparam int TEST_RW1_BYTE_SIZE = 2;
  localparam bit [8:0] TEST_RW1_BYTE_OFFSET = 9'h1f0;
  localparam int TEST_RW1_VAL_BIT_WIDTH = 16;
  localparam bit [15:0] TEST_RW1_VAL_BIT_MASK = 16'hffff;
  localparam int TEST_RW1_VAL_BIT_OFFSET = 0;
  localparam int TEST_RO1_BYTE_WIDTH = 2;
  localparam int TEST_RO1_BYTE_SIZE = 2;
  localparam bit [8:0] TEST_RO1_BYTE_OFFSET = 9'h1f2;
  localparam int TEST_RO1_VAL_BIT_WIDTH = 16;
  localparam bit [15:0] TEST_RO1_VAL_BIT_MASK = 16'hffff;
  localparam int TEST_RO1_VAL_BIT_OFFSET = 0;
  localparam int TEST_RO2_BYTE_WIDTH = 2;
  localparam int TEST_RO2_BYTE_SIZE = 2;
  localparam bit [8:0] TEST_RO2_BYTE_OFFSET = 9'h1f4;
  localparam int TEST_RO2_VAL_BIT_WIDTH = 16;
  localparam bit [15:0] TEST_RO2_VAL_BIT_MASK = 16'hffff;
  localparam int TEST_RO2_VAL_BIT_OFFSET = 0;
  localparam int TEST_RO3_BYTE_WIDTH = 4;
  localparam int TEST_RO3_BYTE_SIZE = 4;
  localparam bit [8:0] TEST_RO3_BYTE_OFFSET = 9'h1f6;
  localparam int TEST_RO3_VAL_BIT_WIDTH = 32;
  localparam bit [31:0] TEST_RO3_VAL_BIT_MASK = 32'hffffffff;
  localparam int TEST_RO3_VAL_BIT_OFFSET = 0;
  localparam int TEST_RO4_BYTE_WIDTH = 4;
  localparam int TEST_RO4_BYTE_SIZE = 4;
  localparam bit [8:0] TEST_RO4_BYTE_OFFSET = 9'h1fa;
  localparam int TEST_RO4_VAL_BIT_WIDTH = 32;
  localparam bit [31:0] TEST_RO4_VAL_BIT_MASK = 32'hffffffff;
  localparam int TEST_RO4_VAL_BIT_OFFSET = 0;
endpackage
