module fastcounter_stage_ #(
    parameter NBITS = 3
) (
    input i_clk,
    input i_rst,
    input i_en,
    input i_load,
    input [NBITS-1:0] i_load_q,
    output [NBITS-1:0] o_q,
    output o_zero
);

    reg [NBITS-1:0] count;
    reg zero;   // registered carry signal

    always @(posedge i_clk or posedge i_rst) begin
        if (i_rst) begin
            count <= {NBITS{1'b0}};
            zero <= 1'b1;
        end else if (i_load) begin
            count <= i_load_q;
            zero <= (i_load_q == {NBITS{1'b0}});
        end else begin
            if (i_en) begin
                count <= count - {{NBITS-1{1'b0}}, 1'b1};
                zero <= (count == {{NBITS-1{1'b0}}, 1'b1});
            end
        end
    end

    assign o_q = count;
    assign o_zero = zero;

endmodule


module fastcounter #(
    parameter NBITS = 10,
    parameter NBITS_STAGE = 9   // default value good for iCE40
) (
    input i_clk,                // clock
    input i_rst,                // assynchronous reset
    //
    input i_en,                 // enable input
    input i_mode,               // mode: 0 - autoreload, 1 - oneshot
    input [NBITS-1:0] i_load_q, // counter load value
    input i_load,               // synchronous counter load (when i_load=1, i_en is ignored)
    //
    output o_zero,              // counter is 0
    output o_nzero,             // counter is not 0
    output o_carry,             // carry pulse
    output o_carry_dly,         // delayed carry pulse
    output o_zpulse,            // zero pulse
    //
    output [NBITS-1:0] o_q      // counter value output
);

    /*****************************************************************************************************************
                        Fast synchronous downcounter

    Fast - because it uses registered carry signals within internal stages, which allows it to obtain
    higher fMAX.

    EN/LOAD/RESET truth table:
         i_rst  i_en  i_load                behavior
           1      *     *       counter loaded with 0, zpulse NOT generated
           0      0     0       no change in state
           0      *     1       counter load: o_q<=i_load_q, zpulse generated if i_load_q==0
           0      1     0       counter decrement (subject to mode and current counter value)

    Modes:
        0 - AUTORELOAD
            if o_q!=0, counter is decremented when i_en==1
            if o_q==0, counter is loaded (o_q<=i_load_q) when i_en==1
        1 - ONESHOT
            if o_q!=0, counter is decremented when i_en==1
            if o_q==0, i_en is disabled, counter may still be reloaded by i_load

    Status outputs:
        o_zero
            is 1 when o_q is zero, 0 otherwise
        o_nzero
            is 1 when o_q is not zero, 0 otherwise
        o_carry
            carry flag
            is 1 when o_q is zero, i_en=1, and counter is not in oneshot mode
        o_carry_dly
            o_carry delayed by 1 i_clk cycle (use to improve timings)
        o_zpulse
            1 clk wide pulse generated when counter value, which was non-zero, becomes zero
            except when counter is reset via i_rst

    Applications:
        In all modes, i_en can be used to "gate" counter decrement. When i_en=0, the counter does not
        decrement (it holds its value unless i_rst or i_load are set), and o_carry is held at 0.
        This can be convenient when counter is driven from another prescaler - in this case, i_en should
        be fed with positive 1x i_clk wide pulses coming at desired count rate.

        Clock prescaler:
            Divides input clock (or frequency of clk gating pulses generated by a different prescaled) by
            DIV_RATIO to generate clk gating pulses with lower frequency.

            i_rst
                Connect to reset network
            i_mode
                set to 0
            i_en
                Divide i_clk: set to 1
                Divide output of another prescaler: connect to output of another prescaler
            i_load
                set to 0
            i_load_q
                set to DIV_RATIO-1, where DIV_RATIO is the desired frequency division ratio
            o_carry, o_carry_dly
                output of prescaler:
                    when DIV_RATIO>1: 1x i_clk wide pulses, one pulse per DIV_RATIO x i_clk or i_en pulses
                    when DIV_RATIO=1: o_carry is a copy of i_en
            o_zero, o_nzero, o_zpulse
                not used

        One-shot:
            When triggered, counter is reloaded with VAL value and then decrements by 1 on each
            i_clk cycle when i_en==1. When counter reaches zero, it stops decrementing till external
            trigger is applied again.

            This allows to generate pulses of specified width, and to generate 1 i_clk wide pulses
            with controlled delay w.r.t trigger.

            Trigger signal is internally processed to make trigger pulse 1x i_clk cycle wide.
            Therefore, increasing trigger pulse width does not cause counter to retrigger or stall.

            i_rst
                Connect to reset network
            i_mode
                set to 1
            i_en
                Count with i_clk rate: set to 1
                Count with prescaled rate: connect to output of prescaler
            i_load
                Connect to positive trigger signal
            i_load_q
                set to NCOUNT
            o_nzero
                Produces positive pulse that starts on the next i_clk cycle after i_load==1
                and has width of NCOUNT i_clk cycles (i_en==1) or i_en pulses (i_en!=1)
            o_zero
                Produces inverted pulse, otherwise same as o_nzero
            o_zpulse
                Produces pulse that is delayed w.r.t. cycle of i_load==1 by NCOUNT+1
                count clocks
            o_carry, o_carry_dly
                not used

    *****************************************************************************************************************/


    localparam MODE_AUTORELOAD = 1'd0;
    localparam MODE_ONESHOT = 1'd1;

    localparam NSTAGES = ((NBITS + NBITS_STAGE - 1) / NBITS_STAGE); // ceil
    localparam NLBITS = NBITS - (NSTAGES-1) * NBITS_STAGE;

    genvar ii;

    // ZERO outputs of all stages
    wire [NSTAGES-1:0] st_zero;
    // EN inputs of all stages
    wire [NSTAGES-1:0] st_en;

    // Shaped load pulse for oneshot mode
    reg load_dly;
    always @(posedge i_clk or posedge i_rst)
        if (i_rst)
            load_dly <= 1'b0;
        else
            load_dly <= i_load;

    wire load_1clk;
    assign load_1clk = i_load && !load_dly;

    // Carry chain logic
    assign st_en[0] = en;
    generate
        for (ii = 1; ii < NSTAGES; ii=ii+1) begin
            assign st_en[ii] = st_zero[ii-1] && st_en[ii-1];
        end
    endgenerate

    // Carry output logic
    assign o_carry = st_en[NSTAGES-1] && st_zero[NSTAGES-1];

    // Delayed carry generator
    reg carry_dly;
    always @(posedge i_clk or posedge i_rst)
        if (i_rst)
            carry_dly <= 1'b0;
        else
            carry_dly <= o_carry;

    assign o_carry_dly = carry_dly;

    // Zero logic
    assign o_zero = & st_zero;    // all stages should be zero
    assign o_nzero = ~o_zero;

    // Mode-dependent enable and load logic
    reg en, load;
    always @(*) begin
        case(i_mode)
        MODE_AUTORELOAD: begin
            en = i_en;
            load = i_load || o_carry;
        end
        default: begin
            // Oneshot
            en = i_en && !o_zero;
            load = load_1clk;
        end
        endcase
    end

    // zpulse generator
    reg zero_dly;
    always @(posedge i_clk or posedge i_rst) begin
        if (i_rst) begin
            zero_dly <= 1'b1;
        end else if (load) begin
            zero_dly <= 1'b0;
        end else begin
            zero_dly <= o_zero;
        end
    end

    assign o_zpulse = o_zero && !zero_dly;

    // Counter stages
    generate
        for (ii = 0; ii < NSTAGES; ii = ii + 1) begin
            if (ii < NSTAGES-1) begin
                fastcounter_stage_ #(
                    .NBITS(NBITS_STAGE)
                ) ctr (
                    .i_clk(i_clk),
                    .i_rst(i_rst),
                    .i_en(st_en[ii]),
                    .i_load(load),
                    .i_load_q(i_load_q[(ii+1)*NBITS_STAGE-1:ii*NBITS_STAGE]),
                    .o_q(o_q[(ii+1)*NBITS_STAGE-1:ii*NBITS_STAGE]),
                    .o_zero(st_zero[ii])
                );
            end else begin
                fastcounter_stage_ #(
                    .NBITS(NLBITS)
                ) ctr (
                    .i_clk(i_clk),
                    .i_rst(i_rst),
                    .i_en(st_en[ii]),
                    .i_load(load),
                    .i_load_q(i_load_q[NBITS-1:ii*NBITS_STAGE]),
                    .o_q(o_q[NBITS-1:ii*NBITS_STAGE]),
                    .o_zero(st_zero[ii])
                );
            end
        end
    endgenerate

endmodule
