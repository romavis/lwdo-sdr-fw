`ifndef LWDO_REGS_VH
`define LWDO_REGS_VH
`define LWDO_REGS_SYS_MAGIC_MAGIC_BIT_WIDTH 32
`define LWDO_REGS_SYS_MAGIC_MAGIC_BIT_MASK 32'hffffffff
`define LWDO_REGS_SYS_MAGIC_MAGIC_BIT_OFFSET 0
`define LWDO_REGS_SYS_MAGIC_BYTE_WIDTH 4
`define LWDO_REGS_SYS_MAGIC_BYTE_SIZE 4
`define LWDO_REGS_SYS_MAGIC_BYTE_OFFSET 9'h000
`define LWDO_REGS_SYS_VERSION_MAJOR_BIT_WIDTH 16
`define LWDO_REGS_SYS_VERSION_MAJOR_BIT_MASK 16'hffff
`define LWDO_REGS_SYS_VERSION_MAJOR_BIT_OFFSET 0
`define LWDO_REGS_SYS_VERSION_MINOR_BIT_WIDTH 16
`define LWDO_REGS_SYS_VERSION_MINOR_BIT_MASK 16'hffff
`define LWDO_REGS_SYS_VERSION_MINOR_BIT_OFFSET 16
`define LWDO_REGS_SYS_VERSION_BYTE_WIDTH 4
`define LWDO_REGS_SYS_VERSION_BYTE_SIZE 4
`define LWDO_REGS_SYS_VERSION_BYTE_OFFSET 9'h004
`define LWDO_REGS_SYS_CON_SYS_RST_BIT_WIDTH 1
`define LWDO_REGS_SYS_CON_SYS_RST_BIT_MASK 1'h1
`define LWDO_REGS_SYS_CON_SYS_RST_BIT_OFFSET 0
`define LWDO_REGS_SYS_CON_BYTE_WIDTH 2
`define LWDO_REGS_SYS_CON_BYTE_SIZE 2
`define LWDO_REGS_SYS_CON_BYTE_OFFSET 9'h008
`define LWDO_REGS_SYS_PLL_DIVR_BIT_WIDTH 4
`define LWDO_REGS_SYS_PLL_DIVR_BIT_MASK 4'hf
`define LWDO_REGS_SYS_PLL_DIVR_BIT_OFFSET 0
`define LWDO_REGS_SYS_PLL_DIVF_BIT_WIDTH 7
`define LWDO_REGS_SYS_PLL_DIVF_BIT_MASK 7'h7f
`define LWDO_REGS_SYS_PLL_DIVF_BIT_OFFSET 4
`define LWDO_REGS_SYS_PLL_DIVQ_BIT_WIDTH 3
`define LWDO_REGS_SYS_PLL_DIVQ_BIT_MASK 3'h7
`define LWDO_REGS_SYS_PLL_DIVQ_BIT_OFFSET 11
`define LWDO_REGS_SYS_PLL_BYTE_WIDTH 2
`define LWDO_REGS_SYS_PLL_BYTE_SIZE 2
`define LWDO_REGS_SYS_PLL_BYTE_OFFSET 9'h00a
`define LWDO_REGS_PDET_CON_EN_BIT_WIDTH 1
`define LWDO_REGS_PDET_CON_EN_BIT_MASK 1'h1
`define LWDO_REGS_PDET_CON_EN_BIT_OFFSET 0
`define LWDO_REGS_PDET_CON_ECLK2_SLOW_BIT_WIDTH 1
`define LWDO_REGS_PDET_CON_ECLK2_SLOW_BIT_MASK 1'h1
`define LWDO_REGS_PDET_CON_ECLK2_SLOW_BIT_OFFSET 1
`define LWDO_REGS_PDET_CON_BYTE_WIDTH 2
`define LWDO_REGS_PDET_CON_BYTE_SIZE 2
`define LWDO_REGS_PDET_CON_BYTE_OFFSET 9'h020
`define LWDO_REGS_PDET_N1_VAL_BIT_WIDTH 32
`define LWDO_REGS_PDET_N1_VAL_BIT_MASK 32'hffffffff
`define LWDO_REGS_PDET_N1_VAL_BIT_OFFSET 0
`define LWDO_REGS_PDET_N1_BYTE_WIDTH 4
`define LWDO_REGS_PDET_N1_BYTE_SIZE 4
`define LWDO_REGS_PDET_N1_BYTE_OFFSET 9'h022
`define LWDO_REGS_PDET_N2_VAL_BIT_WIDTH 32
`define LWDO_REGS_PDET_N2_VAL_BIT_MASK 32'hffffffff
`define LWDO_REGS_PDET_N2_VAL_BIT_OFFSET 0
`define LWDO_REGS_PDET_N2_BYTE_WIDTH 4
`define LWDO_REGS_PDET_N2_BYTE_SIZE 4
`define LWDO_REGS_PDET_N2_BYTE_OFFSET 9'h026
`define LWDO_REGS_ADCT_CON_SRATE1_EN_BIT_WIDTH 1
`define LWDO_REGS_ADCT_CON_SRATE1_EN_BIT_MASK 1'h1
`define LWDO_REGS_ADCT_CON_SRATE1_EN_BIT_OFFSET 0
`define LWDO_REGS_ADCT_CON_SRATE2_EN_BIT_WIDTH 1
`define LWDO_REGS_ADCT_CON_SRATE2_EN_BIT_MASK 1'h1
`define LWDO_REGS_ADCT_CON_SRATE2_EN_BIT_OFFSET 1
`define LWDO_REGS_ADCT_CON_PULS1_EN_BIT_WIDTH 1
`define LWDO_REGS_ADCT_CON_PULS1_EN_BIT_MASK 1'h1
`define LWDO_REGS_ADCT_CON_PULS1_EN_BIT_OFFSET 2
`define LWDO_REGS_ADCT_CON_PULS2_EN_BIT_WIDTH 1
`define LWDO_REGS_ADCT_CON_PULS2_EN_BIT_MASK 1'h1
`define LWDO_REGS_ADCT_CON_PULS2_EN_BIT_OFFSET 3
`define LWDO_REGS_ADCT_CON_BYTE_WIDTH 2
`define LWDO_REGS_ADCT_CON_BYTE_SIZE 2
`define LWDO_REGS_ADCT_CON_BYTE_OFFSET 9'h040
`define LWDO_REGS_ADCT_SRATE1_PSC_DIV_VAL_BIT_WIDTH 8
`define LWDO_REGS_ADCT_SRATE1_PSC_DIV_VAL_BIT_MASK 8'hff
`define LWDO_REGS_ADCT_SRATE1_PSC_DIV_VAL_BIT_OFFSET 0
`define LWDO_REGS_ADCT_SRATE1_PSC_DIV_BYTE_WIDTH 2
`define LWDO_REGS_ADCT_SRATE1_PSC_DIV_BYTE_SIZE 2
`define LWDO_REGS_ADCT_SRATE1_PSC_DIV_BYTE_OFFSET 9'h042
`define LWDO_REGS_ADCT_SRATE2_PSC_DIV_VAL_BIT_WIDTH 8
`define LWDO_REGS_ADCT_SRATE2_PSC_DIV_VAL_BIT_MASK 8'hff
`define LWDO_REGS_ADCT_SRATE2_PSC_DIV_VAL_BIT_OFFSET 0
`define LWDO_REGS_ADCT_SRATE2_PSC_DIV_BYTE_WIDTH 2
`define LWDO_REGS_ADCT_SRATE2_PSC_DIV_BYTE_SIZE 2
`define LWDO_REGS_ADCT_SRATE2_PSC_DIV_BYTE_OFFSET 9'h044
`define LWDO_REGS_ADCT_PULS1_PSC_DIV_VAL_BIT_WIDTH 23
`define LWDO_REGS_ADCT_PULS1_PSC_DIV_VAL_BIT_MASK 23'h7fffff
`define LWDO_REGS_ADCT_PULS1_PSC_DIV_VAL_BIT_OFFSET 0
`define LWDO_REGS_ADCT_PULS1_PSC_DIV_BYTE_WIDTH 4
`define LWDO_REGS_ADCT_PULS1_PSC_DIV_BYTE_SIZE 4
`define LWDO_REGS_ADCT_PULS1_PSC_DIV_BYTE_OFFSET 9'h046
`define LWDO_REGS_ADCT_PULS2_PSC_DIV_VAL_BIT_WIDTH 23
`define LWDO_REGS_ADCT_PULS2_PSC_DIV_VAL_BIT_MASK 23'h7fffff
`define LWDO_REGS_ADCT_PULS2_PSC_DIV_VAL_BIT_OFFSET 0
`define LWDO_REGS_ADCT_PULS2_PSC_DIV_BYTE_WIDTH 4
`define LWDO_REGS_ADCT_PULS2_PSC_DIV_BYTE_SIZE 4
`define LWDO_REGS_ADCT_PULS2_PSC_DIV_BYTE_OFFSET 9'h04a
`define LWDO_REGS_ADCT_PULS1_DLY_VAL_BIT_WIDTH 9
`define LWDO_REGS_ADCT_PULS1_DLY_VAL_BIT_MASK 9'h1ff
`define LWDO_REGS_ADCT_PULS1_DLY_VAL_BIT_OFFSET 0
`define LWDO_REGS_ADCT_PULS1_DLY_BYTE_WIDTH 2
`define LWDO_REGS_ADCT_PULS1_DLY_BYTE_SIZE 2
`define LWDO_REGS_ADCT_PULS1_DLY_BYTE_OFFSET 9'h04e
`define LWDO_REGS_ADCT_PULS2_DLY_VAL_BIT_WIDTH 9
`define LWDO_REGS_ADCT_PULS2_DLY_VAL_BIT_MASK 9'h1ff
`define LWDO_REGS_ADCT_PULS2_DLY_VAL_BIT_OFFSET 0
`define LWDO_REGS_ADCT_PULS2_DLY_BYTE_WIDTH 2
`define LWDO_REGS_ADCT_PULS2_DLY_BYTE_SIZE 2
`define LWDO_REGS_ADCT_PULS2_DLY_BYTE_OFFSET 9'h050
`define LWDO_REGS_ADCT_PULS1_PWIDTH_VAL_BIT_WIDTH 16
`define LWDO_REGS_ADCT_PULS1_PWIDTH_VAL_BIT_MASK 16'hffff
`define LWDO_REGS_ADCT_PULS1_PWIDTH_VAL_BIT_OFFSET 0
`define LWDO_REGS_ADCT_PULS1_PWIDTH_BYTE_WIDTH 2
`define LWDO_REGS_ADCT_PULS1_PWIDTH_BYTE_SIZE 2
`define LWDO_REGS_ADCT_PULS1_PWIDTH_BYTE_OFFSET 9'h052
`define LWDO_REGS_ADCT_PULS2_PWIDTH_VAL_BIT_WIDTH 16
`define LWDO_REGS_ADCT_PULS2_PWIDTH_VAL_BIT_MASK 16'hffff
`define LWDO_REGS_ADCT_PULS2_PWIDTH_VAL_BIT_OFFSET 0
`define LWDO_REGS_ADCT_PULS2_PWIDTH_BYTE_WIDTH 2
`define LWDO_REGS_ADCT_PULS2_PWIDTH_BYTE_SIZE 2
`define LWDO_REGS_ADCT_PULS2_PWIDTH_BYTE_OFFSET 9'h054
`define LWDO_REGS_ADC_CON_ADC1_EN_BIT_WIDTH 1
`define LWDO_REGS_ADC_CON_ADC1_EN_BIT_MASK 1'h1
`define LWDO_REGS_ADC_CON_ADC1_EN_BIT_OFFSET 0
`define LWDO_REGS_ADC_CON_ADC2_EN_BIT_WIDTH 1
`define LWDO_REGS_ADC_CON_ADC2_EN_BIT_MASK 1'h1
`define LWDO_REGS_ADC_CON_ADC2_EN_BIT_OFFSET 1
`define LWDO_REGS_ADC_CON_BYTE_WIDTH 2
`define LWDO_REGS_ADC_CON_BYTE_SIZE 2
`define LWDO_REGS_ADC_CON_BYTE_OFFSET 9'h080
`define LWDO_REGS_ADC_FIFO1_STS_EMPTY_BIT_WIDTH 1
`define LWDO_REGS_ADC_FIFO1_STS_EMPTY_BIT_MASK 1'h1
`define LWDO_REGS_ADC_FIFO1_STS_EMPTY_BIT_OFFSET 0
`define LWDO_REGS_ADC_FIFO1_STS_FULL_BIT_WIDTH 1
`define LWDO_REGS_ADC_FIFO1_STS_FULL_BIT_MASK 1'h1
`define LWDO_REGS_ADC_FIFO1_STS_FULL_BIT_OFFSET 1
`define LWDO_REGS_ADC_FIFO1_STS_HFULL_BIT_WIDTH 1
`define LWDO_REGS_ADC_FIFO1_STS_HFULL_BIT_MASK 1'h1
`define LWDO_REGS_ADC_FIFO1_STS_HFULL_BIT_OFFSET 2
`define LWDO_REGS_ADC_FIFO1_STS_OVFL_BIT_WIDTH 1
`define LWDO_REGS_ADC_FIFO1_STS_OVFL_BIT_MASK 1'h1
`define LWDO_REGS_ADC_FIFO1_STS_OVFL_BIT_OFFSET 3
`define LWDO_REGS_ADC_FIFO1_STS_UDFL_BIT_WIDTH 1
`define LWDO_REGS_ADC_FIFO1_STS_UDFL_BIT_MASK 1'h1
`define LWDO_REGS_ADC_FIFO1_STS_UDFL_BIT_OFFSET 4
`define LWDO_REGS_ADC_FIFO1_STS_BYTE_WIDTH 2
`define LWDO_REGS_ADC_FIFO1_STS_BYTE_SIZE 2
`define LWDO_REGS_ADC_FIFO1_STS_BYTE_OFFSET 9'h082
`define LWDO_REGS_ADC_FIFO2_STS_EMPTY_BIT_WIDTH 1
`define LWDO_REGS_ADC_FIFO2_STS_EMPTY_BIT_MASK 1'h1
`define LWDO_REGS_ADC_FIFO2_STS_EMPTY_BIT_OFFSET 0
`define LWDO_REGS_ADC_FIFO2_STS_FULL_BIT_WIDTH 1
`define LWDO_REGS_ADC_FIFO2_STS_FULL_BIT_MASK 1'h1
`define LWDO_REGS_ADC_FIFO2_STS_FULL_BIT_OFFSET 1
`define LWDO_REGS_ADC_FIFO2_STS_HFULL_BIT_WIDTH 1
`define LWDO_REGS_ADC_FIFO2_STS_HFULL_BIT_MASK 1'h1
`define LWDO_REGS_ADC_FIFO2_STS_HFULL_BIT_OFFSET 2
`define LWDO_REGS_ADC_FIFO2_STS_OVFL_BIT_WIDTH 1
`define LWDO_REGS_ADC_FIFO2_STS_OVFL_BIT_MASK 1'h1
`define LWDO_REGS_ADC_FIFO2_STS_OVFL_BIT_OFFSET 3
`define LWDO_REGS_ADC_FIFO2_STS_UDFL_BIT_WIDTH 1
`define LWDO_REGS_ADC_FIFO2_STS_UDFL_BIT_MASK 1'h1
`define LWDO_REGS_ADC_FIFO2_STS_UDFL_BIT_OFFSET 4
`define LWDO_REGS_ADC_FIFO2_STS_BYTE_WIDTH 2
`define LWDO_REGS_ADC_FIFO2_STS_BYTE_SIZE 2
`define LWDO_REGS_ADC_FIFO2_STS_BYTE_OFFSET 9'h084
`define LWDO_REGS_FTUN_VTUNE_SET_VAL_BIT_WIDTH 16
`define LWDO_REGS_FTUN_VTUNE_SET_VAL_BIT_MASK 16'hffff
`define LWDO_REGS_FTUN_VTUNE_SET_VAL_BIT_OFFSET 0
`define LWDO_REGS_FTUN_VTUNE_SET_BYTE_WIDTH 2
`define LWDO_REGS_FTUN_VTUNE_SET_BYTE_SIZE 2
`define LWDO_REGS_FTUN_VTUNE_SET_BYTE_OFFSET 9'h0a0
`define LWDO_REGS_TEST_RW1_VAL_BIT_WIDTH 16
`define LWDO_REGS_TEST_RW1_VAL_BIT_MASK 16'hffff
`define LWDO_REGS_TEST_RW1_VAL_BIT_OFFSET 0
`define LWDO_REGS_TEST_RW1_BYTE_WIDTH 2
`define LWDO_REGS_TEST_RW1_BYTE_SIZE 2
`define LWDO_REGS_TEST_RW1_BYTE_OFFSET 9'h1f0
`define LWDO_REGS_TEST_RO1_VAL_BIT_WIDTH 16
`define LWDO_REGS_TEST_RO1_VAL_BIT_MASK 16'hffff
`define LWDO_REGS_TEST_RO1_VAL_BIT_OFFSET 0
`define LWDO_REGS_TEST_RO1_BYTE_WIDTH 2
`define LWDO_REGS_TEST_RO1_BYTE_SIZE 2
`define LWDO_REGS_TEST_RO1_BYTE_OFFSET 9'h1f2
`define LWDO_REGS_TEST_RO2_VAL_BIT_WIDTH 16
`define LWDO_REGS_TEST_RO2_VAL_BIT_MASK 16'hffff
`define LWDO_REGS_TEST_RO2_VAL_BIT_OFFSET 0
`define LWDO_REGS_TEST_RO2_BYTE_WIDTH 2
`define LWDO_REGS_TEST_RO2_BYTE_SIZE 2
`define LWDO_REGS_TEST_RO2_BYTE_OFFSET 9'h1f4
`define LWDO_REGS_TEST_RO3_VAL_BIT_WIDTH 32
`define LWDO_REGS_TEST_RO3_VAL_BIT_MASK 32'hffffffff
`define LWDO_REGS_TEST_RO3_VAL_BIT_OFFSET 0
`define LWDO_REGS_TEST_RO3_BYTE_WIDTH 4
`define LWDO_REGS_TEST_RO3_BYTE_SIZE 4
`define LWDO_REGS_TEST_RO3_BYTE_OFFSET 9'h1f6
`define LWDO_REGS_TEST_RO4_VAL_BIT_WIDTH 32
`define LWDO_REGS_TEST_RO4_VAL_BIT_MASK 32'hffffffff
`define LWDO_REGS_TEST_RO4_VAL_BIT_OFFSET 0
`define LWDO_REGS_TEST_RO4_BYTE_WIDTH 4
`define LWDO_REGS_TEST_RO4_BYTE_SIZE 4
`define LWDO_REGS_TEST_RO4_BYTE_OFFSET 9'h1fa
`endif
